CircuitLogix Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 15 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
445 0 1 200 3
126 71 1920 1040
8  5.000 V
8  5.000 V
3 GND
126 71 1920 1040
9437206 0
0
0
0
0
0
0
31
9 Inverter~
13 759 218 0 2 22
0 5 6
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
8953 0 0
0
0
9 Inverter~
13 758 178 0 2 22
0 4 7
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4441 0 0
0
0
9 Inverter~
13 759 138 0 2 22
0 3 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3618 0 0
0
0
9 Inverter~
13 759 98 0 2 22
0 2 9
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
6153 0 0
0
0
9 3-In AND~
219 1019 353 0 4 22
0 8 7 6 10
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 2 0
1 U
5394 0 0
0
0
9 2-In AND~
219 1019 313 0 3 22
0 9 5 12
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7734 0 0
0
0
8 3-In OR~
219 1080 313 0 4 22
0 11 12 10 13
0
0 0 112 0
4 4075
-14 -24 14 -16
0
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 4 0
1 U
9914 0 0
0
0
9 2-In AND~
219 1018 274 0 3 22
0 9 4 11
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3747 0 0
0
0
9 CC 7-Seg~
183 1141 170 0 18 19
10 13 14 15 16 17 18 19 20 21
1 2 2 2 2 2 2 2 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
0
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3549 0 0
0
0
11 Terminal:A~
94 740 98 0 5 9
0 2 2 2 2 22
11 Terminal:A~
19 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
7931 0 0
0
0
11 Terminal:A~
94 720 138 0 5 9
0 3 3 3 3 23
11 Terminal:A~
20 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
9325 0 0
0
0
11 Terminal:A~
94 700 178 0 5 9
0 4 4 4 4 24
11 Terminal:A~
21 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
8903 0 0
0
0
11 Terminal:A~
94 790 218 0 5 9
0 6 6 6 6 25
11 Terminal:A~
22 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3834 0 0
0
0
11 Terminal:A~
94 700 479 0 5 9
0 4 4 4 4 26
11 Terminal:A~
23 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3363 0 0
0
0
11 Terminal:A~
94 680 218 0 5 9
0 5 5 5 5 27
11 Terminal:A~
24 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
7668 0 0
0
0
11 Terminal:A~
94 680 478 0 5 9
0 5 5 5 5 28
11 Terminal:A~
25 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
4718 0 0
0
0
11 Terminal:A~
94 720 479 0 5 9
0 3 3 3 3 29
11 Terminal:A~
26 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3874 0 0
0
0
11 Terminal:A~
94 740 478 0 5 9
0 2 2 2 2 30
11 Terminal:A~
27 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
6671 0 0
0
0
11 Terminal:A~
94 790 218 0 5 9
0 6 6 6 6 31
11 Terminal:A~
28 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3789 0 0
0
0
11 Terminal:A~
94 790 478 0 5 9
0 6 6 6 6 32
11 Terminal:A~
29 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
4871 0 0
0
0
11 Terminal:A~
94 810 178 0 5 9
0 7 7 7 7 33
11 Terminal:A~
30 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3750 0 0
0
0
11 Terminal:A~
94 830 138 0 5 9
0 8 8 8 8 34
11 Terminal:A~
31 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
8778 0 0
0
0
11 Terminal:A~
94 850 98 0 5 9
0 9 9 9 9 35
11 Terminal:A~
32 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
538 0 0
0
0
11 Terminal:A~
94 830 479 0 5 9
0 8 8 8 8 36
11 Terminal:A~
33 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
6843 0 0
0
0
11 Terminal:A~
94 850 478 0 5 9
0 9 9 9 9 37
11 Terminal:A~
34 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
3136 0 0
0
0
11 Terminal:A~
94 810 478 0 5 9
0 7 7 7 7 38
11 Terminal:A~
35 0 16496 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 T
5950 0 0
0
0
14 Logic Display~
6 626 59 0 1 2
10 3
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5670 0 0
0
0
14 Logic Display~
6 648 59 0 1 2
10 2
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6828 0 0
0
0
14 Logic Display~
6 605 59 0 1 2
10 4
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6735 0 0
0
0
14 Logic Display~
6 584 59 0 1 2
10 5
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8365 0 0
0
0
9 Data Seq~
170 540 139 0 17 18
0 39 40 41 42 5 4 3 2 43
44 14 1 16 3 2 0 257
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
0
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
5 SIP10
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
4132 0 0
0
0
AAAAABACADAEAFAGAHAIAJAKALAMANAOAPBABBBCBDBEBFBGBHBIBJBKBLBMBNBOBPCACBCCCDCECFCG
CHCICJCKCLCMCNCOCPDADBDCDDDEDFDGDHDIDJDKDLDMDNDODPEAEBECEDEEEFEGEHEIEJEKELEMENEO
EPFAFBFCFDFEFFFGFHFIFJFKFLFMFNFOFPGAGBGCGDGEGFGGGHGIGJGKGLGMGNGOGPHAHBHCHDHEHFHG
HHHIHJHKHLHMHNHOHPIAIBICIDIEIFIGIHIIIJIKILIMINIOIPJAJBJCJDJEJFJGJHJIJJJKJLJMJNJO
JPKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPLALBLCLDLELFLGLHLILJLKLLLMLNLOLPMAMBMCMDMEMFMG
MHMIMJMKMLMMMNMOMPNANBNCNDNENFNGNHNINJNKNLNMNNNONPOAOBOCODOEOFOGOHOIOJOKOLOMONOO
OPPAPBPCPDPEPFPGPHPIPJPKPLPMPNPOPP
36
1 0 2 0 0 4096 0 28 0 0 8 2
648 77
648 98
1 0 3 0 0 4096 0 27 0 0 7 2
626 77
626 166
1 0 4 0 0 4096 0 29 0 0 6 2
605 77
605 157
1 0 5 0 0 4096 0 30 0 0 5 2
584 77
584 148
3 5 5 0 0 8192 0 15 31 0 0 3
680 213
680 148
572 148
3 6 4 0 0 8192 0 12 31 0 0 3
700 173
700 157
572 157
2 7 3 0 0 0 0 11 31 0 0 4
715 138
639 138
639 166
572 166
2 8 2 0 0 4096 0 10 31 0 0 4
735 98
648 98
648 175
572 175
3 0 6 0 0 4096 0 5 0 0 22 2
995 362
790 362
2 0 7 0 0 4096 0 5 0 0 18 2
995 353
810 353
1 0 8 0 0 4096 0 5 0 0 17 2
995 344
830 344
2 0 5 0 0 4224 0 6 0 0 26 2
995 322
680 322
2 0 4 0 0 4224 0 8 0 0 28 2
994 283
700 283
1 0 9 0 0 4096 0 6 0 0 16 2
995 304
850 304
1 0 9 0 0 0 0 8 0 0 16 2
994 265
850 265
3 1 9 0 0 4224 0 25 23 0 0 2
850 473
850 103
3 1 8 0 0 4224 0 24 22 0 0 2
830 474
830 143
3 1 7 0 0 4224 0 26 21 0 0 2
810 473
810 183
2 2 7 0 0 0 0 2 21 0 0 2
779 178
805 178
2 2 8 0 0 0 0 3 22 0 0 2
780 138
825 138
2 2 9 0 0 0 0 4 23 0 0 2
780 98
845 98
3 1 6 0 0 4224 0 20 13 0 0 2
790 473
790 223
2 2 6 0 0 0 0 19 1 0 0 2
785 218
780 218
1 3 2 0 0 4224 0 10 18 0 0 2
740 103
740 473
1 3 3 0 0 4224 0 11 17 0 0 2
720 143
720 474
1 3 5 0 0 0 0 15 16 0 0 2
680 223
680 473
4 1 5 0 0 0 0 15 1 0 0 2
685 218
744 218
1 3 4 0 0 0 0 12 14 0 0 2
700 183
700 474
2 2 6 0 0 0 0 13 1 0 0 2
785 218
780 218
1 4 4 0 0 0 0 2 12 0 0 2
743 178
705 178
1 4 3 0 0 0 0 3 11 0 0 2
744 138
725 138
1 4 2 0 0 0 0 4 10 0 0 4
744 98
749 98
749 98
745 98
3 4 10 0 0 8320 0 7 5 0 0 4
1067 322
1050 322
1050 353
1040 353
1 3 11 0 0 8320 0 7 8 0 0 4
1067 304
1050 304
1050 274
1039 274
2 3 12 0 0 4224 0 7 6 0 0 2
1068 313
1040 313
1 4 13 0 0 4224 0 9 7 0 0 3
1120 206
1120 313
1113 313
17
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
698 195 713 217
702 199 711 215
1 A
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
698 155 713 177
702 159 711 175
1 B
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
697 116 713 138
701 120 711 136
1 C
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
699 75 715 97
703 79 713 95
1 D
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
637 25 653 47
641 29 651 45
1 D
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
615 25 631 47
621 29 631 45
1 C
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
594 25 609 47
600 29 609 45
1 B
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
574 25 589 47
580 29 589 45
1 A
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
782 480 795 502
786 484 793 500
1 d
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
803 479 816 501
807 483 814 499
1 c
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
821 479 834 501
825 483 832 499
1 b
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
842 478 855 500
846 482 853 498
1 a
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
669 479 685 501
673 483 683 499
1 D
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
690 479 706 501
694 483 704 499
1 C
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
709 479 724 501
713 483 722 499
1 B
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 1
729 479 744 501
733 483 742 499
1 A
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 27
1037 94 1219 116
1043 98 1219 114
27 Vicent van Gogh - CG3015678
0
0 2 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.032 5e-006 5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
