CircuitLogix Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1263 30 100 3
126 71 1366 720
7 5.000 V
7 5.000 V
3 GND
126 71 1366 720
9437202 0
0
0
0
0
0
0
96
13 Logic Switch~
5 242 1428 0 1 3
0 12
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 240 1402 0 1 3
0 9
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 243 1367 0 1 3
0 7
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3618 0 0
0
0
13 Logic Switch~
5 241 1340 0 1 3
0 88
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -2 0
1 V
6153 0 0
0
0
13 Logic Switch~
5 240 1174 0 1 3
0 22
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5394 0 0
0
0
13 Logic Switch~
5 238 1148 0 1 3
0 23
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7734 0 0
0
0
13 Logic Switch~
5 241 1113 0 1 3
0 24
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9914 0 0
0
0
13 Logic Switch~
5 239 1086 0 1 3
0 28
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3747 0 0
0
0
13 Logic Switch~
5 234 923 0 1 3
0 34
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3549 0 0
0
0
13 Logic Switch~
5 232 897 0 1 3
0 38
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7931 0 0
0
0
13 Logic Switch~
5 235 862 0 1 3
0 36
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9325 0 0
0
0
13 Logic Switch~
5 233 835 0 1 3
0 33
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8903 0 0
0
0
13 Logic Switch~
5 238 738 0 1 3
0 53
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3834 0 0
0
0
13 Logic Switch~
5 236 712 0 1 3
0 50
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3363 0 0
0
0
13 Logic Switch~
5 239 677 0 1 3
0 56
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7668 0 0
0
0
13 Logic Switch~
5 237 650 0 1 3
0 48
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4718 0 0
0
0
13 Logic Switch~
5 229 548 0 1 3
0 63
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3874 0 0
0
0
13 Logic Switch~
5 227 522 0 1 3
0 64
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6671 0 0
0
0
13 Logic Switch~
5 230 487 0 1 3
0 67
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3789 0 0
0
0
13 Logic Switch~
5 228 460 0 1 3
0 65
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4871 0 0
0
0
13 Logic Switch~
5 215 227 0 1 3
0 75
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3750 0 0
0
0
13 Logic Switch~
5 213 201 0 1 3
0 76
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8778 0 0
0
0
13 Logic Switch~
5 216 166 0 1 3
0 77
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
538 0 0
0
0
13 Logic Switch~
5 214 139 0 1 3
0 78
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6843 0 0
0
0
13 Logic Switch~
5 220 396 0 1 3
0 81
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3136 0 0
0
0
13 Logic Switch~
5 218 370 0 1 3
0 87
0
0 0 20848 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5950 0 0
0
0
13 Logic Switch~
5 221 335 0 1 3
0 85
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5670 0 0
0
0
13 Logic Switch~
5 219 308 0 1 3
0 89
0
0 0 20848 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 0 0 -1 0
1 V
6828 0 0
0
0
14 Logic Display~
6 520 1390 0 1 2
10 2
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6735 0 0
0
0
9 Inverter~
13 477 1424 0 2 22
0 6 2
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 22 0
1 U
8365 0 0
0
0
9 3-In NOR~
219 413 1425 0 4 22
0 5 4 3 6
0
0 0 112 0
6 74LS27
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 11 10 9 8 0
65 0 0 0 3 2 20 0
1 U
4132 0 0
0
0
9 Inverter~
13 280 1365 0 2 22
0 7 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 22 0
1 U
4551 0 0
0
0
9 2-In AND~
219 341 1376 0 3 22
0 8 9 5
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
3635 0 0
0
0
9 Inverter~
13 287 1479 0 2 22
0 9 10
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 22 0
1 U
3973 0 0
0
0
9 Inverter~
13 282 1454 0 2 22
0 9 11
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
3851 0 0
0
0
9 2-In AND~
219 343 1465 0 3 22
0 11 10 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
8383 0 0
0
0
9 2-In AND~
219 344 1420 0 3 22
0 9 12 4
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
9334 0 0
0
0
9 Inverter~
13 9 1075 0 2 22
0 90 91
0
0 0 112 90
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 512 6 6 19 0
1 U
7471 0 0
0
0
14 Logic Display~
6 590 1135 0 1 2
10 13
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3334 0 0
0
0
8 2-In OR~
219 534 1159 0 3 22
0 15 14 13
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
3559 0 0
0
0
8 2-In OR~
219 429 1232 0 3 22
0 18 17 14
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
984 0 0
0
0
9 Inverter~
13 497 1109 0 2 22
0 16 15
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 19 0
1 U
7557 0 0
0
0
9 3-In NOR~
219 433 1110 0 4 22
0 21 20 19 16
0
0 0 112 0
6 74LS27
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 11 10 9 8 0
65 0 0 0 3 1 20 0
1 U
3146 0 0
0
0
9 Inverter~
13 338 1286 0 2 22
0 22 26
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 19 0
1 U
5687 0 0
0
0
9 Inverter~
13 332 1256 0 2 22
0 23 25
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 19 0
1 U
7939 0 0
0
0
5 7415~
219 381 1256 0 4 22
0 24 25 26 17
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 18 0
1 U
3308 0 0
0
0
9 2-In AND~
219 374 1207 0 3 22
0 23 22 18
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
3408 0 0
0
0
9 Inverter~
13 278 1120 0 2 22
0 24 27
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 13 0
1 U
9773 0 0
0
0
9 2-In AND~
219 376 1163 0 3 22
0 27 22 19
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
691 0 0
0
0
9 2-In AND~
219 376 1121 0 3 22
0 28 22 20
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
7834 0 0
0
0
9 Inverter~
13 271 1087 0 2 22
0 28 29
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 13 0
1 U
3588 0 0
0
0
9 2-In AND~
219 361 1086 0 3 22
0 29 23 21
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
4528 0 0
0
0
5 7415~
219 387 892 0 4 22
0 33 32 31 30
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 15 0
1 U
3303 0 0
0
0
9 Inverter~
13 284 916 0 2 22
0 34 31
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 13 0
1 U
9654 0 0
0
0
14 Logic Display~
6 628 901 0 1 2
10 39
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9791 0 0
0
0
8 2-In OR~
219 574 930 0 3 22
0 41 40 39
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
4589 0 0
0
0
9 Inverter~
13 521 891 0 2 22
0 44 41
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 13 0
1 U
964 0 0
0
0
9 3-In NOR~
219 460 891 0 4 22
0 43 30 42 44
0
0 0 112 0
6 74LS27
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 10 9 8 1 2 13 12 3
4 5 6 11 10 9 8 0
65 0 0 0 3 3 10 0
1 U
9151 0 0
0
0
8 2-In OR~
219 470 1011 0 3 22
0 46 45 40
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
4745 0 0
0
0
5 7415~
219 404 1029 0 4 22
0 33 35 34 45
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 15 0
1 U
8433 0 0
0
0
5 7415~
219 405 983 0 4 22
0 37 38 31 46
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 15 0
1 U
4221 0 0
0
0
9 4-In AND~
219 400 946 0 5 22
0 37 36 32 31 42
0
0 0 112 0
6 74LS21
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 1 14 0
1 U
8348 0 0
0
0
9 Inverter~
13 288 884 0 2 22
0 38 32
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
5299 0 0
0
0
9 Inverter~
13 285 856 0 2 22
0 36 35
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
7393 0 0
0
0
9 Inverter~
13 285 833 0 2 22
0 33 37
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
6917 0 0
0
0
9 4-In AND~
219 406 841 0 5 22
0 37 35 32 34 43
0
0 0 112 0
6 74LS21
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 2 11 0
1 U
8767 0 0
0
0
14 Logic Display~
6 577 638 0 1 2
10 47
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3606 0 0
0
0
9 2-In AND~
219 423 656 0 3 22
0 48 50 49
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6970 0 0
0
0
5 7415~
219 437 734 0 4 22
0 54 50 53 52
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 2 7 0
1 U
343 0 0
0
0
9 Inverter~
13 302 775 0 2 22
0 53 57
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
7197 0 0
0
0
9 Inverter~
13 297 730 0 2 22
0 50 58
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3623 0 0
0
0
9 Inverter~
13 294 701 0 2 22
0 56 54
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
7656 0 0
0
0
9 Inverter~
13 296 675 0 2 22
0 48 59
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
5365 0 0
0
0
9 4-In AND~
219 386 704 0 5 22
0 59 54 58 57 55
0
0 0 112 0
6 74LS21
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 -961104021
65 0 0 0 2 1 11 0
1 U
4557 0 0
0
0
9 Inverter~
13 550 688 0 2 22
0 51 47
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
3489 0 0
0
0
9 3-In NOR~
219 495 687 0 4 22
0 49 55 52 51
0
0 0 112 0
6 74LS27
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 4 5 6 1 2 13 12 3
4 5 6 11 10 9 8 0
65 0 0 0 3 2 10 0
1 U
345 0 0
0
0
14 Logic Display~
6 577 475 0 1 2
10 60
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3374 0 0
0
0
9 4-In AND~
219 422 550 0 5 22
0 65 66 64 63 61
0
0 0 112 0
6 74LS21
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 -961104021
65 0 0 0 2 2 3 0
1 U
5866 0 0
0
0
9 Inverter~
13 303 559 0 2 22
0 67 66
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
631 0 0
0
0
9 Inverter~
13 291 524 0 2 22
0 64 68
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
745 0 0
0
0
9 2-In AND~
219 386 519 0 3 22
0 65 68 62
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
7222 0 0
0
0
9 Inverter~
13 527 489 0 2 22
0 70 60
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
4508 0 0
0
0
9 3-In NOR~
219 461 489 0 4 22
0 69 62 61 70
0
0 0 112 0
6 74LS27
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 11 10 9 8 0
65 0 0 0 3 1 10 0
1 U
3738 0 0
0
0
9 3-In AND~
219 372 479 0 4 22
0 71 64 63 69
0
0 0 112 0
6 74LS11
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 9 0
1 U
91 0 0
0
0
9 Inverter~
13 273 463 0 2 22
0 65 71
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
4965 0 0
0
0
14 Logic Display~
6 502 122 0 1 2
10 72
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7791 0 0
0
0
9 4-In AND~
219 365 136 0 5 22
0 78 77 76 75 74
0
0 0 112 0
6 74LS21
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
16

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0
65 0 0 0 2 1 3 0
1 U
3467 0 0
0
0
8 2-In OR~
219 432 153 0 3 22
0 74 73 72
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3907 0 0
0
0
5 7415~
219 369 190 0 4 22
0 77 76 79 73
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 1 7 0
1 U
7505 0 0
0
0
9 Inverter~
13 270 227 0 2 22
0 75 79
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 4 0
1 U
6423 0 0
0
0
9 Inverter~
13 283 400 0 2 22
0 81 80
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 4 0
1 U
3623 0 0
0
0
14 Logic Display~
6 498 339 0 1 2
10 82
0
0 0 53344 0
6 100MEG
10 -16 38 -8
0
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8523 0 0
0
0
5 7415~
219 367 385 0 4 22
0 85 86 80 83
0
0 0 112 0
6 74LS15
-21 -28 21 -20
0
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0
65 0 0 0 3 3 5 0
1 U
9623 0 0
0
0
9 Inverter~
13 285 376 0 2 22
0 87 86
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 4 0
1 U
9468 0 0
0
0
8 2-In OR~
219 454 366 0 3 22
0 84 83 82
0
0 0 112 0
6 74LS32
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
9254 0 0
0
0
9 2-In AND~
219 380 344 0 3 22
0 85 81 84
0
0 0 112 0
6 74LS08
-21 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5587 0 0
0
0
124
1 2 2 0 0 8320 0 29 30 0 0 3
520 1408
520 1424
498 1424
3 3 3 0 0 8320 0 31 36 0 0 4
400 1434
372 1434
372 1465
364 1465
2 3 4 0 0 4224 0 31 37 0 0 4
401 1425
373 1425
373 1420
365 1420
1 3 5 0 0 8320 0 31 33 0 0 4
400 1416
370 1416
370 1376
362 1376
1 4 6 0 0 8320 0 30 31 0 0 3
462 1424
462 1425
452 1425
1 1 7 0 0 8320 0 32 3 0 0 3
265 1365
265 1367
255 1367
1 2 8 0 0 4224 0 33 32 0 0 4
317 1367
309 1367
309 1365
301 1365
2 0 9 0 0 4096 0 33 0 0 9 4
317 1385
266 1385
266 1402
261 1402
1 0 9 0 0 8320 0 34 0 0 11 3
272 1479
261 1479
261 1402
2 2 10 0 0 12416 0 36 34 0 0 4
319 1474
316 1474
316 1479
308 1479
1 0 9 0 0 0 0 35 0 0 14 5
267 1454
261 1454
261 1438
260 1438
261 1402
1 2 11 0 0 4224 0 36 35 0 0 4
319 1456
310 1456
310 1454
303 1454
2 1 12 0 0 4224 0 37 1 0 0 4
320 1429
263 1429
263 1428
254 1428
1 1 9 0 0 0 0 37 2 0 0 4
320 1411
261 1411
261 1402
252 1402
3 1 13 0 0 4224 0 40 39 0 0 3
567 1159
590 1159
590 1153
3 2 14 0 0 8320 0 41 40 0 0 4
462 1232
513 1232
513 1168
521 1168
2 1 15 0 0 8320 0 42 40 0 0 6
518 1109
522 1109
522 1140
516 1140
516 1150
521 1150
1 4 16 0 0 8320 0 42 43 0 0 3
482 1109
482 1110
472 1110
2 4 17 0 0 8320 0 41 46 0 0 4
416 1241
410 1241
410 1256
402 1256
1 3 18 0 0 8320 0 41 47 0 0 4
416 1223
403 1223
403 1207
395 1207
3 3 19 0 0 8320 0 43 49 0 0 4
420 1119
405 1119
405 1163
397 1163
2 3 20 0 0 4224 0 43 50 0 0 4
421 1110
405 1110
405 1121
397 1121
1 3 21 0 0 4224 0 43 52 0 0 4
420 1101
390 1101
390 1086
382 1086
1 1 22 0 0 8320 0 44 5 0 0 4
323 1286
261 1286
261 1174
252 1174
1 0 23 0 0 8320 0 45 0 0 36 3
317 1256
291 1256
291 1148
1 1 24 0 0 4224 0 46 7 0 0 3
357 1247
357 1113
253 1113
2 2 25 0 0 4224 0 45 46 0 0 2
353 1256
357 1256
2 3 26 0 0 4224 0 44 46 0 0 3
359 1286
359 1265
357 1265
2 0 22 0 0 0 0 47 0 0 31 4
350 1216
268 1216
268 1174
263 1174
1 0 23 0 0 0 0 47 0 0 36 3
350 1198
279 1198
279 1148
2 0 22 0 0 0 0 49 0 0 34 4
352 1172
352 1181
263 1181
263 1174
1 1 24 0 0 0 0 48 7 0 0 3
263 1120
263 1113
253 1113
1 2 27 0 0 4224 0 49 48 0 0 4
352 1154
312 1154
312 1120
299 1120
2 1 22 0 0 0 0 50 5 0 0 3
352 1130
352 1174
252 1174
1 1 28 0 0 8320 0 50 8 0 0 4
352 1112
352 1106
251 1106
251 1086
1 2 23 0 0 0 0 6 52 0 0 4
250 1148
305 1148
305 1095
337 1095
1 1 28 0 0 0 0 51 8 0 0 3
256 1087
256 1086
251 1086
2 1 29 0 0 12416 0 51 52 0 0 4
292 1087
305 1087
305 1077
337 1077
4 2 30 0 0 4224 0 53 58 0 0 4
408 892
439 892
439 891
448 891
3 2 31 0 0 4096 0 53 54 0 0 4
363 901
313 901
313 916
305 916
2 2 32 0 0 4096 0 53 63 0 0 4
363 892
317 892
317 884
309 884
1 0 33 0 0 8192 0 53 0 0 45 3
363 883
363 858
260 858
3 0 34 0 0 8320 0 60 0 0 53 4
380 1038
264 1038
264 919
266 919
2 2 35 0 0 8320 0 60 64 0 0 4
380 1029
314 1029
314 856
306 856
1 0 33 0 0 8320 0 60 0 0 54 3
380 1020
260 1020
260 833
3 2 31 0 0 8320 0 61 54 0 0 4
381 992
313 992
313 916
305 916
4 2 31 0 0 0 0 62 54 0 0 4
376 960
313 960
313 916
305 916
3 2 32 0 0 8320 0 62 63 0 0 4
376 951
317 951
317 884
309 884
2 0 36 0 0 4224 0 62 0 0 55 3
376 942
258 942
258 856
1 0 37 0 0 8192 0 62 0 0 60 5
376 933
314 933
314 833
306 833
306 828
2 0 38 0 0 4224 0 61 0 0 56 3
381 983
258 983
258 884
1 0 37 0 0 8320 0 61 0 0 60 3
381 974
314 974
314 828
1 0 34 0 0 0 0 54 0 0 57 4
269 916
266 917
266 923
255 923
1 1 33 0 0 0 0 65 12 0 0 4
270 833
257 833
257 835
245 835
1 1 36 0 0 0 0 64 11 0 0 4
270 856
256 856
256 862
247 862
1 1 38 0 0 0 0 63 10 0 0 4
273 884
253 884
253 897
244 897
4 1 34 0 0 0 0 66 9 0 0 6
382 855
336 855
336 937
255 937
255 923
246 923
3 2 32 0 0 0 0 66 63 0 0 4
382 846
326 846
326 884
309 884
2 2 35 0 0 0 0 66 64 0 0 4
382 837
318 837
318 856
306 856
1 2 37 0 0 0 0 66 65 0 0 3
382 828
306 828
306 833
3 1 39 0 0 4224 0 56 55 0 0 3
607 930
628 930
628 919
2 3 40 0 0 8320 0 56 59 0 0 4
561 939
511 939
511 1011
503 1011
1 2 41 0 0 8320 0 56 57 0 0 4
561 921
544 921
544 891
542 891
3 5 42 0 0 8320 0 58 62 0 0 4
447 900
438 900
438 946
421 946
1 5 43 0 0 8320 0 58 66 0 0 4
447 882
438 882
438 841
427 841
4 1 44 0 0 4224 0 58 57 0 0 4
499 891
507 891
507 891
506 891
2 4 45 0 0 4224 0 59 60 0 0 4
457 1020
433 1020
433 1029
425 1029
1 4 46 0 0 4224 0 59 61 0 0 4
457 1002
436 1002
436 983
426 983
1 2 47 0 0 4224 0 67 75 0 0 3
577 656
577 688
571 688
1 0 48 0 0 4224 0 68 0 0 82 4
399 647
273 647
273 660
258 660
3 1 49 0 0 8320 0 68 76 0 0 3
444 656
444 678
482 678
2 0 50 0 0 4224 0 68 0 0 80 4
399 665
262 665
262 723
257 723
4 1 51 0 0 4224 0 76 75 0 0 4
534 687
538 687
538 688
535 688
4 3 52 0 0 8320 0 69 76 0 0 6
458 734
462 734
462 703
453 703
453 696
482 696
3 0 53 0 0 8320 0 69 0 0 79 3
413 743
413 757
259 757
2 0 50 0 0 0 0 69 0 0 80 4
413 734
322 734
322 715
257 715
1 2 54 0 0 8320 0 69 72 0 0 3
413 725
413 701
315 701
5 2 55 0 0 4224 0 74 76 0 0 4
407 704
450 704
450 687
483 687
1 1 53 0 0 0 0 70 13 0 0 4
287 775
259 775
259 738
250 738
1 1 50 0 0 0 0 71 14 0 0 4
282 730
257 730
257 712
248 712
1 1 56 0 0 8320 0 72 15 0 0 4
279 701
260 701
260 677
251 677
1 1 48 0 0 0 0 73 16 0 0 4
281 675
258 675
258 650
249 650
2 4 57 0 0 8320 0 70 74 0 0 4
323 775
354 775
354 718
362 718
2 3 58 0 0 4224 0 71 74 0 0 4
318 730
354 730
354 709
362 709
2 2 54 0 0 0 0 72 74 0 0 5
315 701
315 703
354 703
354 700
362 700
2 1 59 0 0 4224 0 73 74 0 0 4
317 675
354 675
354 691
362 691
2 1 60 0 0 4224 0 82 77 0 0 5
548 489
565 489
565 490
577 490
577 493
5 3 61 0 0 8320 0 78 83 0 0 6
443 550
447 550
447 508
443 508
443 498
448 498
2 3 62 0 0 4224 0 83 81 0 0 4
449 489
415 489
415 519
407 519
4 1 63 0 0 12288 0 78 17 0 0 6
398 564
328 564
328 544
250 544
250 548
241 548
3 1 64 0 0 12288 0 78 18 0 0 6
398 555
328 555
328 509
248 509
248 522
239 522
1 1 65 0 0 12416 0 78 20 0 0 6
398 537
411 537
411 448
249 448
249 460
240 460
2 2 66 0 0 4224 0 79 78 0 0 4
324 559
429 559
429 546
398 546
1 1 67 0 0 8320 0 79 19 0 0 4
288 559
251 559
251 487
242 487
1 0 65 0 0 0 0 81 0 0 103 3
362 510
251 510
251 463
2 2 68 0 0 4224 0 80 81 0 0 4
312 524
354 524
354 528
362 528
1 1 64 0 0 0 0 80 18 0 0 4
276 524
248 524
248 522
239 522
4 1 69 0 0 4224 0 84 83 0 0 4
393 479
440 479
440 480
448 480
1 4 70 0 0 4224 0 82 83 0 0 2
512 489
500 489
3 1 63 0 0 4224 0 84 17 0 0 4
348 488
250 488
250 548
241 548
2 1 64 0 0 4224 0 84 18 0 0 4
348 479
248 479
248 522
239 522
2 1 71 0 0 4224 0 85 84 0 0 4
294 463
344 463
344 470
348 470
1 1 65 0 0 0 0 85 20 0 0 4
258 463
249 463
249 460
240 460
1 3 72 0 0 8320 0 86 88 0 0 3
502 140
502 153
465 153
4 2 73 0 0 8320 0 89 88 0 0 4
390 190
411 190
411 162
419 162
5 1 74 0 0 4224 0 87 88 0 0 4
386 136
411 136
411 144
419 144
4 1 75 0 0 4224 0 87 21 0 0 4
341 150
236 150
236 227
227 227
3 1 76 0 0 4096 0 87 22 0 0 4
341 141
234 141
234 201
225 201
2 1 77 0 0 4096 0 87 23 0 0 4
341 132
237 132
237 166
228 166
1 1 78 0 0 4224 0 24 87 0 0 4
226 139
333 139
333 123
341 123
1 1 75 0 0 0 0 90 21 0 0 2
255 227
227 227
3 2 79 0 0 4224 0 89 90 0 0 4
345 199
299 199
299 227
291 227
2 1 76 0 0 4224 0 89 22 0 0 4
345 190
234 190
234 201
225 201
1 1 77 0 0 4224 0 89 23 0 0 4
345 181
237 181
237 166
228 166
2 3 80 0 0 4224 0 91 93 0 0 4
304 400
335 400
335 394
343 394
1 0 81 0 0 4096 0 91 0 0 123 4
268 400
246 400
246 388
241 388
1 3 82 0 0 8320 0 92 95 0 0 3
498 357
498 366
487 366
4 2 83 0 0 4224 0 93 95 0 0 4
388 385
433 385
433 375
441 375
3 1 84 0 0 4224 0 96 95 0 0 4
401 344
433 344
433 357
441 357
1 0 85 0 0 8192 0 93 0 0 124 3
343 376
343 339
259 339
2 2 86 0 0 4224 0 94 93 0 0 4
306 376
335 376
335 385
343 385
1 1 87 0 0 4224 0 26 94 0 0 4
230 370
262 370
262 376
270 376
2 1 81 0 0 4224 0 96 25 0 0 4
356 353
241 353
241 396
232 396
1 1 85 0 0 4224 0 96 27 0 0 6
356 335
259 335
259 339
232 339
232 335
233 335
6
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 2
595 1128 611 1150
606 1136 616 1152
2 sf
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 2
647 888 667 910
658 896 672 912
2 se
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 2
586 629 606 651
597 637 611 653
2 sd
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 2
593 469 613 491
604 477 618 493
2 sc
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 2
502 114 522 136
513 122 527 138
2 sa
16 6 0 0 0 0 0 0 0 0 0 0 39
5 Arial
0 0 0 3
494 336 516 358
505 343 521 359
3 sb'
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
